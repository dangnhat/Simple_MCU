library verilog;
use verilog.vl_types.all;
entity testbench_CPU is
end testbench_CPU;
